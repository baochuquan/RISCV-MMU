library verilog;
use verilog.vl_types.all;
entity PTW is
    generic(
        S_ready         : vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi0);
        S_req           : vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi1);
        S_wait1         : vl_logic_vector(0 to 2) := (Hi0, Hi1, Hi0);
        S_wait2         : vl_logic_vector(0 to 2) := (Hi0, Hi1, Hi1);
        S_set_dirty     : vl_logic_vector(0 to 2) := (Hi1, Hi0, Hi0);
        S_wait1_dirty   : vl_logic_vector(0 to 2) := (Hi1, Hi0, Hi1);
        S_wait2_dirty   : vl_logic_vector(0 to 2) := (Hi1, Hi1, Hi0);
        S_done          : vl_logic_vector(0 to 2) := (Hi1, Hi1, Hi1)
    );
    port(
        clock           : in     vl_logic;
        reset           : in     vl_logic;
        io_requestor_0_req_ready: out    vl_logic;
        io_requestor_0_req_valid: in     vl_logic;
        io_requestor_0_req_bits_prv: in     vl_logic_vector(1 downto 0);
        io_requestor_0_req_bits_pum: in     vl_logic;
        io_requestor_0_req_bits_mxr: in     vl_logic;
        io_requestor_0_req_bits_addr: in     vl_logic_vector(26 downto 0);
        io_requestor_0_req_bits_store: in     vl_logic;
        io_requestor_0_req_bits_fetch: in     vl_logic;
        io_requestor_0_resp_valid: out    vl_logic;
        io_requestor_0_resp_bits_pte_reserved_for_hardware: out    vl_logic_vector(15 downto 0);
        io_requestor_0_resp_bits_pte_ppn: out    vl_logic_vector(37 downto 0);
        io_requestor_0_resp_bits_pte_reserved_for_software: out    vl_logic_vector(1 downto 0);
        io_requestor_0_resp_bits_pte_d: out    vl_logic;
        io_requestor_0_resp_bits_pte_a: out    vl_logic;
        io_requestor_0_resp_bits_pte_g: out    vl_logic;
        io_requestor_0_resp_bits_pte_u: out    vl_logic;
        io_requestor_0_resp_bits_pte_x: out    vl_logic;
        io_requestor_0_resp_bits_pte_w: out    vl_logic;
        io_requestor_0_resp_bits_pte_r: out    vl_logic;
        io_requestor_0_resp_bits_pte_v: out    vl_logic;
        io_requestor_0_ptbr_asid: out    vl_logic_vector(6 downto 0);
        io_requestor_0_ptbr_ppn: out    vl_logic_vector(37 downto 0);
        io_requestor_0_invalidate: out    vl_logic;
        io_requestor_0_status_debug: out    vl_logic;
        io_requestor_0_status_isa: out    vl_logic_vector(31 downto 0);
        io_requestor_0_status_prv: out    vl_logic_vector(1 downto 0);
        io_requestor_0_status_sd: out    vl_logic;
        io_requestor_0_status_zero3: out    vl_logic_vector(30 downto 0);
        io_requestor_0_status_sd_rv32: out    vl_logic;
        io_requestor_0_status_zero2: out    vl_logic_vector(1 downto 0);
        io_requestor_0_status_vm: out    vl_logic_vector(4 downto 0);
        io_requestor_0_status_zero1: out    vl_logic_vector(3 downto 0);
        io_requestor_0_status_mxr: out    vl_logic;
        io_requestor_0_status_pum: out    vl_logic;
        io_requestor_0_status_mprv: out    vl_logic;
        io_requestor_0_status_xs: out    vl_logic_vector(1 downto 0);
        io_requestor_0_status_fs: out    vl_logic_vector(1 downto 0);
        io_requestor_0_status_mpp: out    vl_logic_vector(1 downto 0);
        io_requestor_0_status_hpp: out    vl_logic_vector(1 downto 0);
        io_requestor_0_status_spp: out    vl_logic;
        io_requestor_0_status_mpie: out    vl_logic;
        io_requestor_0_status_hpie: out    vl_logic;
        io_requestor_0_status_spie: out    vl_logic;
        io_requestor_0_status_upie: out    vl_logic;
        io_requestor_0_status_mie: out    vl_logic;
        io_requestor_0_status_hie: out    vl_logic;
        io_requestor_0_status_sie: out    vl_logic;
        io_requestor_0_status_uie: out    vl_logic;
        io_requestor_1_req_ready: out    vl_logic;
        io_requestor_1_req_valid: in     vl_logic;
        io_requestor_1_req_bits_prv: in     vl_logic_vector(1 downto 0);
        io_requestor_1_req_bits_pum: in     vl_logic;
        io_requestor_1_req_bits_mxr: in     vl_logic;
        io_requestor_1_req_bits_addr: in     vl_logic_vector(26 downto 0);
        io_requestor_1_req_bits_store: in     vl_logic;
        io_requestor_1_req_bits_fetch: in     vl_logic;
        io_requestor_1_resp_valid: out    vl_logic;
        io_requestor_1_resp_bits_pte_reserved_for_hardware: out    vl_logic_vector(15 downto 0);
        io_requestor_1_resp_bits_pte_ppn: out    vl_logic_vector(37 downto 0);
        io_requestor_1_resp_bits_pte_reserved_for_software: out    vl_logic_vector(1 downto 0);
        io_requestor_1_resp_bits_pte_d: out    vl_logic;
        io_requestor_1_resp_bits_pte_a: out    vl_logic;
        io_requestor_1_resp_bits_pte_g: out    vl_logic;
        io_requestor_1_resp_bits_pte_u: out    vl_logic;
        io_requestor_1_resp_bits_pte_x: out    vl_logic;
        io_requestor_1_resp_bits_pte_w: out    vl_logic;
        io_requestor_1_resp_bits_pte_r: out    vl_logic;
        io_requestor_1_resp_bits_pte_v: out    vl_logic;
        io_requestor_1_ptbr_asid: out    vl_logic_vector(6 downto 0);
        io_requestor_1_ptbr_ppn: out    vl_logic_vector(37 downto 0);
        io_requestor_1_invalidate: out    vl_logic;
        io_requestor_1_status_debug: out    vl_logic;
        io_requestor_1_status_isa: out    vl_logic_vector(31 downto 0);
        io_requestor_1_status_prv: out    vl_logic_vector(1 downto 0);
        io_requestor_1_status_sd: out    vl_logic;
        io_requestor_1_status_zero3: out    vl_logic_vector(30 downto 0);
        io_requestor_1_status_sd_rv32: out    vl_logic;
        io_requestor_1_status_zero2: out    vl_logic_vector(1 downto 0);
        io_requestor_1_status_vm: out    vl_logic_vector(4 downto 0);
        io_requestor_1_status_zero1: out    vl_logic_vector(3 downto 0);
        io_requestor_1_status_mxr: out    vl_logic;
        io_requestor_1_status_pum: out    vl_logic;
        io_requestor_1_status_mprv: out    vl_logic;
        io_requestor_1_status_xs: out    vl_logic_vector(1 downto 0);
        io_requestor_1_status_fs: out    vl_logic_vector(1 downto 0);
        io_requestor_1_status_mpp: out    vl_logic_vector(1 downto 0);
        io_requestor_1_status_hpp: out    vl_logic_vector(1 downto 0);
        io_requestor_1_status_spp: out    vl_logic;
        io_requestor_1_status_mpie: out    vl_logic;
        io_requestor_1_status_hpie: out    vl_logic;
        io_requestor_1_status_spie: out    vl_logic;
        io_requestor_1_status_upie: out    vl_logic;
        io_requestor_1_status_mie: out    vl_logic;
        io_requestor_1_status_hie: out    vl_logic;
        io_requestor_1_status_sie: out    vl_logic;
        io_requestor_1_status_uie: out    vl_logic;
        io_mem_req_ready: in     vl_logic;
        io_mem_req_valid: out    vl_logic;
        io_mem_req_bits_addr: out    vl_logic_vector(39 downto 0);
        io_mem_req_bits_tag: out    vl_logic_vector(6 downto 0);
        io_mem_req_bits_cmd: out    vl_logic_vector(4 downto 0);
        io_mem_req_bits_typ: out    vl_logic_vector(2 downto 0);
        io_mem_req_bits_phys: out    vl_logic;
        io_mem_req_bits_data: out    vl_logic_vector(63 downto 0);
        io_mem_s1_kill  : out    vl_logic;
        io_mem_s1_data  : out    vl_logic_vector(63 downto 0);
        io_mem_s2_nack  : in     vl_logic;
        io_mem_resp_valid: in     vl_logic;
        io_mem_resp_bits_data: in     vl_logic_vector(63 downto 0);
        io_mem_xcpt_pf_ld: in     vl_logic;
        io_mem_xcpt_pf_st: in     vl_logic;
        io_mem_invalidate_lr: out    vl_logic;
        io_mem_ordered  : in     vl_logic;
        io_dpath_ptbr_asid: in     vl_logic_vector(6 downto 0);
        io_dpath_ptbr_ppn: in     vl_logic_vector(37 downto 0);
        io_dpath_invalidate: in     vl_logic;
        io_dpath_status_debug: in     vl_logic;
        io_dpath_status_isa: in     vl_logic_vector(31 downto 0);
        io_dpath_status_prv: in     vl_logic_vector(1 downto 0);
        io_dpath_status_sd: in     vl_logic;
        io_dpath_status_zero3: in     vl_logic_vector(30 downto 0);
        io_dpath_status_sd_rv32: in     vl_logic;
        io_dpath_status_zero2: in     vl_logic_vector(1 downto 0);
        io_dpath_status_vm: in     vl_logic_vector(4 downto 0);
        io_dpath_status_zero1: in     vl_logic_vector(3 downto 0);
        io_dpath_status_mxr: in     vl_logic;
        io_dpath_status_pum: in     vl_logic;
        io_dpath_status_mprv: in     vl_logic;
        io_dpath_status_xs: in     vl_logic_vector(1 downto 0);
        io_dpath_status_fs: in     vl_logic_vector(1 downto 0);
        io_dpath_status_mpp: in     vl_logic_vector(1 downto 0);
        io_dpath_status_hpp: in     vl_logic_vector(1 downto 0);
        io_dpath_status_spp: in     vl_logic;
        io_dpath_status_mpie: in     vl_logic;
        io_dpath_status_hpie: in     vl_logic;
        io_dpath_status_spie: in     vl_logic;
        io_dpath_status_upie: in     vl_logic;
        io_dpath_status_mie: in     vl_logic;
        io_dpath_status_hie: in     vl_logic;
        io_dpath_status_sie: in     vl_logic;
        io_dpath_status_uie: in     vl_logic
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of S_ready : constant is 1;
    attribute mti_svvh_generic_type of S_req : constant is 1;
    attribute mti_svvh_generic_type of S_wait1 : constant is 1;
    attribute mti_svvh_generic_type of S_wait2 : constant is 1;
    attribute mti_svvh_generic_type of S_set_dirty : constant is 1;
    attribute mti_svvh_generic_type of S_wait1_dirty : constant is 1;
    attribute mti_svvh_generic_type of S_wait2_dirty : constant is 1;
    attribute mti_svvh_generic_type of S_done : constant is 1;
end PTW;
