module standard_PTW(
  input   clock,
  input   reset,
  output  io_requestor_0_req_ready,
  input   io_requestor_0_req_valid,
  input  [1:0] io_requestor_0_req_bits_prv,
  input   io_requestor_0_req_bits_pum,
  input   io_requestor_0_req_bits_mxr,
  input  [26:0] io_requestor_0_req_bits_addr,
  input   io_requestor_0_req_bits_store,
  input   io_requestor_0_req_bits_fetch,
  output  io_requestor_0_resp_valid,
  output [15:0] io_requestor_0_resp_bits_pte_reserved_for_hardware,
  output [37:0] io_requestor_0_resp_bits_pte_ppn,
  output [1:0] io_requestor_0_resp_bits_pte_reserved_for_software,
  output  io_requestor_0_resp_bits_pte_d,
  output  io_requestor_0_resp_bits_pte_a,
  output  io_requestor_0_resp_bits_pte_g,
  output  io_requestor_0_resp_bits_pte_u,
  output  io_requestor_0_resp_bits_pte_x,
  output  io_requestor_0_resp_bits_pte_w,
  output  io_requestor_0_resp_bits_pte_r,
  output  io_requestor_0_resp_bits_pte_v,
  output [6:0] io_requestor_0_ptbr_asid,
  output [37:0] io_requestor_0_ptbr_ppn,
  output  io_requestor_0_invalidate,
  output  io_requestor_0_status_debug,
  output [31:0] io_requestor_0_status_isa,
  output [1:0] io_requestor_0_status_prv,
  output  io_requestor_0_status_sd,
  output [30:0] io_requestor_0_status_zero3,
  output  io_requestor_0_status_sd_rv32,
  output [1:0] io_requestor_0_status_zero2,
  output [4:0] io_requestor_0_status_vm,
  output [3:0] io_requestor_0_status_zero1,
  output  io_requestor_0_status_mxr,
  output  io_requestor_0_status_pum,
  output  io_requestor_0_status_mprv,
  output [1:0] io_requestor_0_status_xs,
  output [1:0] io_requestor_0_status_fs,
  output [1:0] io_requestor_0_status_mpp,
  output [1:0] io_requestor_0_status_hpp,
  output  io_requestor_0_status_spp,
  output  io_requestor_0_status_mpie,
  output  io_requestor_0_status_hpie,
  output  io_requestor_0_status_spie,
  output  io_requestor_0_status_upie,
  output  io_requestor_0_status_mie,
  output  io_requestor_0_status_hie,
  output  io_requestor_0_status_sie,
  output  io_requestor_0_status_uie,
  output  io_requestor_1_req_ready,
  input   io_requestor_1_req_valid,
  input  [1:0] io_requestor_1_req_bits_prv,
  input   io_requestor_1_req_bits_pum,
  input   io_requestor_1_req_bits_mxr,
  input  [26:0] io_requestor_1_req_bits_addr,
  input   io_requestor_1_req_bits_store,
  input   io_requestor_1_req_bits_fetch,
  output  io_requestor_1_resp_valid,
  output [15:0] io_requestor_1_resp_bits_pte_reserved_for_hardware,
  output [37:0] io_requestor_1_resp_bits_pte_ppn,
  output [1:0] io_requestor_1_resp_bits_pte_reserved_for_software,
  output  io_requestor_1_resp_bits_pte_d,
  output  io_requestor_1_resp_bits_pte_a,
  output  io_requestor_1_resp_bits_pte_g,
  output  io_requestor_1_resp_bits_pte_u,
  output  io_requestor_1_resp_bits_pte_x,
  output  io_requestor_1_resp_bits_pte_w,
  output  io_requestor_1_resp_bits_pte_r,
  output  io_requestor_1_resp_bits_pte_v,
  output [6:0] io_requestor_1_ptbr_asid,
  output [37:0] io_requestor_1_ptbr_ppn,
  output  io_requestor_1_invalidate,
  output  io_requestor_1_status_debug,
  output [31:0] io_requestor_1_status_isa,
  output [1:0] io_requestor_1_status_prv,
  output  io_requestor_1_status_sd,
  output [30:0] io_requestor_1_status_zero3,
  output  io_requestor_1_status_sd_rv32,
  output [1:0] io_requestor_1_status_zero2,
  output [4:0] io_requestor_1_status_vm,
  output [3:0] io_requestor_1_status_zero1,
  output  io_requestor_1_status_mxr,
  output  io_requestor_1_status_pum,
  output  io_requestor_1_status_mprv,
  output [1:0] io_requestor_1_status_xs,
  output [1:0] io_requestor_1_status_fs,
  output [1:0] io_requestor_1_status_mpp,
  output [1:0] io_requestor_1_status_hpp,
  output  io_requestor_1_status_spp,
  output  io_requestor_1_status_mpie,
  output  io_requestor_1_status_hpie,
  output  io_requestor_1_status_spie,
  output  io_requestor_1_status_upie,
  output  io_requestor_1_status_mie,
  output  io_requestor_1_status_hie,
  output  io_requestor_1_status_sie,
  output  io_requestor_1_status_uie,
  input   io_mem_req_ready,
  output  io_mem_req_valid,
  output [39:0] io_mem_req_bits_addr,
  output [6:0] io_mem_req_bits_tag,
  output [4:0] io_mem_req_bits_cmd,
  output [2:0] io_mem_req_bits_typ,
  output  io_mem_req_bits_phys,
  output [63:0] io_mem_req_bits_data,
  output  io_mem_s1_kill,
  output [63:0] io_mem_s1_data,
  input   io_mem_s2_nack,
  input   io_mem_resp_valid,/*
  input  [39:0] io_mem_resp_bits_addr,
  input  [6:0] io_mem_resp_bits_tag,
  input  [4:0] io_mem_resp_bits_cmd,
  input  [2:0] io_mem_resp_bits_typ,*/
  input  [63:0] io_mem_resp_bits_data,/*
  input   io_mem_resp_bits_replay,
  input   io_mem_resp_bits_has_data,
  input  [63:0] io_mem_resp_bits_data_word_bypass,
  input  [63:0] io_mem_resp_bits_store_data,
  input   io_mem_replay_next,
  input   io_mem_xcpt_ma_ld,
  input   io_mem_xcpt_ma_st,*/
  input   io_mem_xcpt_pf_ld,
  input   io_mem_xcpt_pf_st,
  output  io_mem_invalidate_lr,
  input   io_mem_ordered,
  input  [6:0] io_dpath_ptbr_asid,
  input  [37:0] io_dpath_ptbr_ppn,
  input   io_dpath_invalidate,
  input   io_dpath_status_debug,
  input  [31:0] io_dpath_status_isa,
  input  [1:0] io_dpath_status_prv,
  input   io_dpath_status_sd,
  input  [30:0] io_dpath_status_zero3,
  input   io_dpath_status_sd_rv32,
  input  [1:0] io_dpath_status_zero2,
  input  [4:0] io_dpath_status_vm,
  input  [3:0] io_dpath_status_zero1,
  input   io_dpath_status_mxr,
  input   io_dpath_status_pum,
  input   io_dpath_status_mprv,
  input  [1:0] io_dpath_status_xs,
  input  [1:0] io_dpath_status_fs,
  input  [1:0] io_dpath_status_mpp,
  input  [1:0] io_dpath_status_hpp,
  input   io_dpath_status_spp,
  input   io_dpath_status_mpie,
  input   io_dpath_status_hpie,
  input   io_dpath_status_spie,
  input   io_dpath_status_upie,
  input   io_dpath_status_mie,
  input   io_dpath_status_hie,
  input   io_dpath_status_sie,
  input   io_dpath_status_uie
);
  reg [2:0] state;
  reg [31:0] GEN_125;
  reg [1:0] count;
  reg [31:0] GEN_126;
  reg  s1_kill;
  reg [31:0] GEN_127;
  reg [1:0] r_req_prv;
  reg [31:0] GEN_128;
  reg  r_req_pum;
  reg [31:0] GEN_129;
  reg  r_req_mxr;
  reg [31:0] GEN_130;
  reg [26:0] r_req_addr;
  reg [31:0] GEN_131;
  reg  r_req_store;
  reg [31:0] GEN_132;
  reg  r_req_fetch;
  reg [31:0] GEN_133;
  reg  r_req_dest;
  reg [31:0] GEN_134;
  reg [15:0] r_pte_reserved_for_hardware;
  reg [31:0] GEN_135;
  reg [37:0] r_pte_ppn;
  reg [63:0] GEN_136;
  reg [1:0] r_pte_reserved_for_software;
  reg [31:0] GEN_137;
  reg  r_pte_d;
  reg [31:0] GEN_138;
  reg  r_pte_a;
  reg [31:0] GEN_139;
  reg  r_pte_g;
  reg [31:0] GEN_140;
  reg  r_pte_u;
  reg [31:0] GEN_141;
  reg  r_pte_x;
  reg [31:0] GEN_142;
  reg  r_pte_w;
  reg [31:0] GEN_143;
  reg  r_pte_r;
  reg [31:0] GEN_144;
  reg  r_pte_v;
  reg [31:0] GEN_145;
  wire [8:0] T_2207;
  wire [17:0] T_2208;
  wire [8:0] vpn_idxs_1;
  wire [8:0] vpn_idxs_2;
  wire [1:0] T_2211;
  wire  T_2213;
  wire  T_2217;
  wire [8:0] T_2218;
  wire [8:0] vpn_idx;
  wire  arb_clock;
  wire  arb_reset;
  wire  arb_io_in_0_ready;
  wire  arb_io_in_0_valid;
  wire [1:0] arb_io_in_0_bits_prv;
  wire  arb_io_in_0_bits_pum;
  wire  arb_io_in_0_bits_mxr;
  wire [26:0] arb_io_in_0_bits_addr;
  wire  arb_io_in_0_bits_store;
  wire  arb_io_in_0_bits_fetch;
  wire  arb_io_in_1_ready;
  wire  arb_io_in_1_valid;
  wire [1:0] arb_io_in_1_bits_prv;
  wire  arb_io_in_1_bits_pum;
  wire  arb_io_in_1_bits_mxr;
  wire [26:0] arb_io_in_1_bits_addr;
  wire  arb_io_in_1_bits_store;
  wire  arb_io_in_1_bits_fetch;
  wire  arb_io_out_ready;
  wire  arb_io_out_valid;
  wire [1:0] arb_io_out_bits_prv;
  wire  arb_io_out_bits_pum;
  wire  arb_io_out_bits_mxr;
  wire [26:0] arb_io_out_bits_addr;
  wire  arb_io_out_bits_store;
  wire  arb_io_out_bits_fetch;
  wire  arb_io_chosen;
  wire  T_2226;
  wire [15:0] T_2251_reserved_for_hardware;
  wire [37:0] T_2251_ppn;
  wire [1:0] T_2251_reserved_for_software;
  wire  T_2251_d;
  wire  T_2251_a;
  wire  T_2251_g;
  wire  T_2251_u;
  wire  T_2251_x;
  wire  T_2251_w;
  wire  T_2251_r;
  wire  T_2251_v;
  wire  T_2263;
  wire  T_2264;
  wire  T_2265;
  wire  T_2266;
  wire  T_2267;
  wire  T_2268;
  wire  T_2269;
  wire  T_2270;
  wire [1:0] T_2271;
  wire [37:0] T_2272;
  wire [15:0] T_2273;
  wire [15:0] T_2298_reserved_for_hardware;
  wire [37:0] T_2298_ppn;
  wire [1:0] T_2298_reserved_for_software;
  wire  T_2298_d;
  wire  T_2298_a;
  wire  T_2298_g;
  wire  T_2298_u;
  wire  T_2298_x;
  wire  T_2298_w;
  wire  T_2298_r;
  wire  T_2298_v;
  wire [15:0] pte_reserved_for_hardware;
  wire [37:0] pte_ppn;
  wire [1:0] pte_reserved_for_software;
  wire  pte_d;
  wire  pte_a;
  wire  pte_g;
  wire  pte_u;
  wire  pte_x;
  wire  pte_w;
  wire  pte_r;
  wire  pte_v;
  wire [19:0] T_2332;
  wire [17:0] T_2333;
  wire  T_2335;
  wire  GEN_2;
  wire [46:0] T_2337;
  wire [49:0] GEN_113;
  wire [49:0] pte_addr;
  wire  T_2338;
  wire [1:0] GEN_3;
  wire  GEN_4;
  wire  GEN_5;
  wire [26:0] GEN_6;
  wire  GEN_7;
  wire  GEN_8;
  wire  GEN_9;
  wire [37:0] GEN_10;
  reg [7:0] T_2340;
  reg [31:0] GEN_146;
  reg [7:0] T_2342;
  reg [31:0] GEN_147;
  reg [31:0] T_2349_0;
  reg [31:0] GEN_148;
  reg [31:0] T_2349_1;
  reg [31:0] GEN_149;
  reg [31:0] T_2349_2;
  reg [31:0] GEN_150;
  reg [31:0] T_2349_3;
  reg [31:0] GEN_151;
  reg [31:0] T_2349_4;
  reg [31:0] GEN_152;
  reg [31:0] T_2349_5;
  reg [31:0] GEN_153;
  reg [31:0] T_2349_6;
  reg [31:0] GEN_154;
  reg [31:0] T_2349_7;
  reg [31:0] GEN_155;
  reg [19:0] T_2357_0;
  reg [31:0] GEN_156;
  reg [19:0] T_2357_1;
  reg [31:0] GEN_157;
  reg [19:0] T_2357_2;
  reg [31:0] GEN_158;
  reg [19:0] T_2357_3;
  reg [31:0] GEN_159;
  reg [19:0] T_2357_4;
  reg [31:0] GEN_160;
  reg [19:0] T_2357_5;
  reg [31:0] GEN_161;
  reg [19:0] T_2357_6;
  reg [31:0] GEN_162;
  reg [19:0] T_2357_7;
  reg [31:0] GEN_163;
  wire [49:0] GEN_114;
  wire  T_2359;
  wire [49:0] GEN_115;
  wire  T_2360;
  wire [49:0] GEN_116;
  wire  T_2361;
  wire [49:0] GEN_117;
  wire  T_2362;
  wire [49:0] GEN_118;
  wire  T_2363;
  wire [49:0] GEN_119;
  wire  T_2364;
  wire [49:0] GEN_120;
  wire  T_2365;
  wire [49:0] GEN_121;
  wire  T_2366;
  wire [1:0] T_2367;
  wire [1:0] T_2368;
  wire [3:0] T_2369;
  wire [1:0] T_2370;
  wire [1:0] T_2371;
  wire [3:0] T_2372;
  wire [7:0] T_2373;
  wire [7:0] T_2374;
  wire  T_2376;
  wire  T_2378;
  wire  T_2379;
  wire  T_2381;
  wire  T_2382;
  wire  T_2384;
  wire  T_2385;
  wire  T_2386;
  wire  T_2388;
  wire  T_2389;
  wire [7:0] T_2390;
  wire  T_2392;
  wire [7:0] T_2394;
  wire  T_2395;
  wire [1:0] T_2396;
  wire [7:0] T_2397;
  wire  T_2398;
  wire [2:0] T_2399;
  wire [7:0] T_2400;
  wire  T_2401;
  wire [3:0] T_2402;
  wire [2:0] T_2403;
  wire  T_2405;
  wire  T_2406;
  wire  T_2407;
  wire  T_2408;
  wire  T_2409;
  wire  T_2410;
  wire  T_2411;
  wire [2:0] T_2421;
  wire [2:0] T_2422;
  wire [2:0] T_2423;
  wire [2:0] T_2424;
  wire [2:0] T_2425;
  wire [2:0] T_2426;
  wire [2:0] T_2427;
  wire [2:0] T_2428;
  wire [7:0] T_2430;
  wire [7:0] T_2431;
  wire [31:0] GEN_0;
  wire [31:0] GEN_11;
  wire [31:0] GEN_12;
  wire [31:0] GEN_13;
  wire [31:0] GEN_14;
  wire [31:0] GEN_15;
  wire [31:0] GEN_16;
  wire [31:0] GEN_17;
  wire [31:0] GEN_18;
  wire [19:0] GEN_1;
  wire [19:0] GEN_19;
  wire [19:0] GEN_20;
  wire [19:0] GEN_21;
  wire [19:0] GEN_22;
  wire [19:0] GEN_23;
  wire [19:0] GEN_24;
  wire [19:0] GEN_25;
  wire [19:0] GEN_26;
  wire [7:0] GEN_27;
  wire [31:0] GEN_28;
  wire [31:0] GEN_29;
  wire [31:0] GEN_30;
  wire [31:0] GEN_31;
  wire [31:0] GEN_32;
  wire [31:0] GEN_33;
  wire [31:0] GEN_34;
  wire [31:0] GEN_35;
  wire [19:0] GEN_36;
  wire [19:0] GEN_37;
  wire [19:0] GEN_38;
  wire [19:0] GEN_39;
  wire [19:0] GEN_40;
  wire [19:0] GEN_41;
  wire [19:0] GEN_42;
  wire [19:0] GEN_43;
  wire  T_2432;
  wire  T_2433;
  wire [3:0] T_2434;
  wire [3:0] T_2435;
  wire  T_2437;
  wire [3:0] T_2438;
  wire [1:0] T_2439;
  wire [1:0] T_2440;
  wire  T_2442;
  wire [1:0] T_2443;
  wire  T_2444;
  wire [1:0] T_2445;
  wire [2:0] T_2446;
  wire  T_2448;
  wire  T_2450;
  wire [1:0] T_2452;
  wire [7:0] GEN_122;
  wire [7:0] T_2453;
  wire [7:0] T_2454;
  wire [7:0] T_2455;
  wire [7:0] T_2456;
  wire [7:0] T_2457;
  wire [1:0] T_2458;
  wire  T_2459;
  wire  T_2461;
  wire [3:0] T_2463;
  wire [7:0] GEN_124;
  wire [7:0] T_2464;
  wire [7:0] T_2465;
  wire [7:0] T_2466;
  wire [7:0] T_2467;
  wire [7:0] T_2468;
  wire [2:0] T_2469;
  wire  T_2470;
  wire  T_2472;
  wire [7:0] T_2474;
  wire [7:0] T_2475;
  wire [7:0] T_2476;
  wire [7:0] T_2477;
  wire [7:0] T_2478;
  wire [7:0] T_2479;
  wire [7:0] GEN_44;
  wire [7:0] GEN_45;
  wire  T_2483;
  wire  pte_cache_hit;
  wire  T_2484;
  wire  T_2485;
  wire  T_2486;
  wire  T_2487;
  wire  T_2488;
  wire  T_2489;
  wire  T_2490;
  wire  T_2491;
  wire [19:0] T_2493;
  wire [19:0] T_2495;
  wire [19:0] T_2497;
  wire [19:0] T_2499;
  wire [19:0] T_2501;
  wire [19:0] T_2503;
  wire [19:0] T_2505;
  wire [19:0] T_2507;
  wire [19:0] T_2509;
  wire [19:0] T_2510;
  wire [19:0] T_2511;
  wire [19:0] T_2512;
  wire [19:0] T_2513;
  wire [19:0] T_2514;
  wire [19:0] T_2515;
  wire [19:0] pte_cache_data;
  wire [15:0] T_2541_reserved_for_hardware;
  wire [37:0] T_2541_ppn;
  wire [1:0] T_2541_reserved_for_software;
  wire  T_2541_d;
  wire  T_2541_a;
  wire  T_2541_g;
  wire  T_2541_u;
  wire  T_2541_x;
  wire  T_2541_w;
  wire  T_2541_r;
  wire  T_2541_v;
  wire [63:0] T_2554;
  wire  T_2555;
  wire  T_2556;
  wire  T_2557;
  wire  T_2558;
  wire  T_2559;
  wire  T_2560;
  wire  T_2561;
  wire  T_2562;
  wire [1:0] T_2563;
  wire [37:0] T_2564;
  wire [15:0] T_2565;
  wire [15:0] pte_wdata_reserved_for_hardware;
  wire [37:0] pte_wdata_ppn;
  wire [1:0] pte_wdata_reserved_for_software;
  wire  pte_wdata_d;
  wire  pte_wdata_a;
  wire  pte_wdata_g;
  wire  pte_wdata_u;
  wire  pte_wdata_x;
  wire  pte_wdata_w;
  wire  pte_wdata_r;
  wire  pte_wdata_v;
  wire  T_2579;
  wire  T_2580;
  wire [4:0] T_2583;
  wire [1:0] T_2585;
  wire [1:0] T_2586;
  wire [2:0] T_2587;
  wire [4:0] T_2588;
  wire [1:0] T_2589;
  wire [2:0] T_2590;
  wire [53:0] T_2591;
  wire [55:0] T_2592;
  wire [58:0] T_2593;
  wire [63:0] T_2594;
  wire [19:0] T_2596;
  wire [17:0] T_2597;
  wire [37:0] resp_ppns_0;
  wire [28:0] T_2598;
  wire [37:0] resp_ppns_1;
  wire [37:0] resp_ppns_2;
  wire  T_2600;
  wire  T_2602;
  wire  T_2603;
  wire [37:0] T_2612;
  wire [37:0] T_2613;
  wire  T_2617;
  wire  T_2628;
  wire [2:0] GEN_46;
  wire [2:0] GEN_47;
  wire [1:0] GEN_48;
  wire  T_2630;
  wire [2:0] T_2633;
  wire [1:0] T_2634;
  wire [2:0] GEN_50;
  wire [1:0] GEN_51;
  wire [37:0] GEN_52;
  wire  T_2636;
  wire  T_2637;
  wire [2:0] GEN_53;
  wire  GEN_54;
  wire [2:0] GEN_55;
  wire [1:0] GEN_56;
  wire [37:0] GEN_57;
  wire  T_2638;
  wire  GEN_58;
  wire [2:0] GEN_59;
  wire [2:0] GEN_60;
  wire  GEN_61;
  wire  T_2640;
  wire [2:0] GEN_62;
  wire  T_2641;
  wire  T_2642;
  wire  T_2643;
  wire  T_2644;
  wire  T_2646;
  wire  T_2647;
  wire  T_2648;
  wire  T_2651;
  wire  T_2652;
  wire  T_2653;
  wire  T_2654;
  wire  T_2655;
  wire  T_2657;
  wire  T_2659;
  wire  T_2660;
  wire  T_2661;
  wire  T_2662;
  wire [2:0] GEN_63;
  wire  T_2664;
  wire [15:0] GEN_64;
  wire [37:0] GEN_65;
  wire [1:0] GEN_66;
  wire  GEN_67;
  wire  GEN_68;
  wire  GEN_69;
  wire  GEN_70;
  wire  GEN_71;
  wire  GEN_72;
  wire  GEN_73;
  wire  GEN_74;
  wire  T_2676;
  wire [2:0] GEN_75;
  wire [1:0] GEN_76;
  wire [2:0] GEN_77;
  wire [15:0] GEN_78;
  wire [37:0] GEN_79;
  wire [1:0] GEN_80;
  wire  GEN_81;
  wire  GEN_82;
  wire  GEN_83;
  wire  GEN_84;
  wire  GEN_85;
  wire  GEN_86;
  wire  GEN_87;
  wire  GEN_88;
  wire [1:0] GEN_89;
  wire [2:0] GEN_90;
  wire [15:0] GEN_91;
  wire [37:0] GEN_92;
  wire [1:0] GEN_93;
  wire  GEN_94;
  wire  GEN_95;
  wire  GEN_96;
  wire  GEN_97;
  wire  GEN_98;
  wire  GEN_99;
  wire  GEN_100;
  wire  GEN_101;
  wire [1:0] GEN_102;
  wire  T_2680;
  wire [2:0] GEN_103;
  wire [2:0] GEN_104;
  wire  T_2681;
  wire  GEN_105;
  wire [2:0] GEN_106;
  wire [2:0] GEN_107;
  wire  GEN_108;
  wire  T_2683;
  wire [2:0] GEN_109;
  wire [2:0] GEN_110;
  wire [2:0] GEN_111;
  wire  T_2684;
  wire [2:0] GEN_112;
  reg [6:0] GEN_49;
  reg [31:0] GEN_164;
  reg [63:0] GEN_123;
  reg [63:0] GEN_165;
  RRArbiter arb (
    .clock(arb_clock),
    .reset(arb_reset),
    .io_in_0_ready(arb_io_in_0_ready),
    .io_in_0_valid(arb_io_in_0_valid),
    .io_in_0_bits_prv(arb_io_in_0_bits_prv),
    .io_in_0_bits_pum(arb_io_in_0_bits_pum),
    .io_in_0_bits_mxr(arb_io_in_0_bits_mxr),
    .io_in_0_bits_addr(arb_io_in_0_bits_addr),
    .io_in_0_bits_store(arb_io_in_0_bits_store),
    .io_in_0_bits_fetch(arb_io_in_0_bits_fetch),
    .io_in_1_ready(arb_io_in_1_ready),
    .io_in_1_valid(arb_io_in_1_valid),
    .io_in_1_bits_prv(arb_io_in_1_bits_prv),
    .io_in_1_bits_pum(arb_io_in_1_bits_pum),
    .io_in_1_bits_mxr(arb_io_in_1_bits_mxr),
    .io_in_1_bits_addr(arb_io_in_1_bits_addr),
    .io_in_1_bits_store(arb_io_in_1_bits_store),
    .io_in_1_bits_fetch(arb_io_in_1_bits_fetch),
    .io_out_ready(arb_io_out_ready),
    .io_out_valid(arb_io_out_valid),
    .io_out_bits_prv(arb_io_out_bits_prv),
    .io_out_bits_pum(arb_io_out_bits_pum),
    .io_out_bits_mxr(arb_io_out_bits_mxr),
    .io_out_bits_addr(arb_io_out_bits_addr),
    .io_out_bits_store(arb_io_out_bits_store),
    .io_out_bits_fetch(arb_io_out_bits_fetch),
    .io_chosen(arb_io_chosen)
  );
  assign io_requestor_0_req_ready = arb_io_in_0_ready;
  assign io_requestor_0_resp_valid = T_2603;
  assign io_requestor_0_resp_bits_pte_reserved_for_hardware = r_pte_reserved_for_hardware;
  assign io_requestor_0_resp_bits_pte_ppn = T_2613;
  assign io_requestor_0_resp_bits_pte_reserved_for_software = r_pte_reserved_for_software;
  assign io_requestor_0_resp_bits_pte_d = r_pte_d;
  assign io_requestor_0_resp_bits_pte_a = r_pte_a;
  assign io_requestor_0_resp_bits_pte_g = r_pte_g;
  assign io_requestor_0_resp_bits_pte_u = r_pte_u;
  assign io_requestor_0_resp_bits_pte_x = r_pte_x;
  assign io_requestor_0_resp_bits_pte_w = r_pte_w;
  assign io_requestor_0_resp_bits_pte_r = r_pte_r;
  assign io_requestor_0_resp_bits_pte_v = r_pte_v;
  assign io_requestor_0_ptbr_asid = io_dpath_ptbr_asid;
  assign io_requestor_0_ptbr_ppn = io_dpath_ptbr_ppn;
  assign io_requestor_0_invalidate = io_dpath_invalidate;
  assign io_requestor_0_status_debug = io_dpath_status_debug;
  assign io_requestor_0_status_isa = io_dpath_status_isa;
  assign io_requestor_0_status_prv = io_dpath_status_prv;
  assign io_requestor_0_status_sd = io_dpath_status_sd;
  assign io_requestor_0_status_zero3 = io_dpath_status_zero3;
  assign io_requestor_0_status_sd_rv32 = io_dpath_status_sd_rv32;
  assign io_requestor_0_status_zero2 = io_dpath_status_zero2;
  assign io_requestor_0_status_vm = io_dpath_status_vm;
  assign io_requestor_0_status_zero1 = io_dpath_status_zero1;
  assign io_requestor_0_status_mxr = io_dpath_status_mxr;
  assign io_requestor_0_status_pum = io_dpath_status_pum;
  assign io_requestor_0_status_mprv = io_dpath_status_mprv;
  assign io_requestor_0_status_xs = io_dpath_status_xs;
  assign io_requestor_0_status_fs = io_dpath_status_fs;
  assign io_requestor_0_status_mpp = io_dpath_status_mpp;
  assign io_requestor_0_status_hpp = io_dpath_status_hpp;
  assign io_requestor_0_status_spp = io_dpath_status_spp;
  assign io_requestor_0_status_mpie = io_dpath_status_mpie;
  assign io_requestor_0_status_hpie = io_dpath_status_hpie;
  assign io_requestor_0_status_spie = io_dpath_status_spie;
  assign io_requestor_0_status_upie = io_dpath_status_upie;
  assign io_requestor_0_status_mie = io_dpath_status_mie;
  assign io_requestor_0_status_hie = io_dpath_status_hie;
  assign io_requestor_0_status_sie = io_dpath_status_sie;
  assign io_requestor_0_status_uie = io_dpath_status_uie;
  assign io_requestor_1_req_ready = arb_io_in_1_ready;
  assign io_requestor_1_resp_valid = T_2617;
  assign io_requestor_1_resp_bits_pte_reserved_for_hardware = r_pte_reserved_for_hardware;
  assign io_requestor_1_resp_bits_pte_ppn = T_2613;
  assign io_requestor_1_resp_bits_pte_reserved_for_software = r_pte_reserved_for_software;
  assign io_requestor_1_resp_bits_pte_d = r_pte_d;
  assign io_requestor_1_resp_bits_pte_a = r_pte_a;
  assign io_requestor_1_resp_bits_pte_g = r_pte_g;
  assign io_requestor_1_resp_bits_pte_u = r_pte_u;
  assign io_requestor_1_resp_bits_pte_x = r_pte_x;
  assign io_requestor_1_resp_bits_pte_w = r_pte_w;
  assign io_requestor_1_resp_bits_pte_r = r_pte_r;
  assign io_requestor_1_resp_bits_pte_v = r_pte_v;
  assign io_requestor_1_ptbr_asid = io_dpath_ptbr_asid;
  assign io_requestor_1_ptbr_ppn = io_dpath_ptbr_ppn;
  assign io_requestor_1_invalidate = io_dpath_invalidate;
  assign io_requestor_1_status_debug = io_dpath_status_debug;
  assign io_requestor_1_status_isa = io_dpath_status_isa;
  assign io_requestor_1_status_prv = io_dpath_status_prv;
  assign io_requestor_1_status_sd = io_dpath_status_sd;
  assign io_requestor_1_status_zero3 = io_dpath_status_zero3;
  assign io_requestor_1_status_sd_rv32 = io_dpath_status_sd_rv32;
  assign io_requestor_1_status_zero2 = io_dpath_status_zero2;
  assign io_requestor_1_status_vm = io_dpath_status_vm;
  assign io_requestor_1_status_zero1 = io_dpath_status_zero1;
  assign io_requestor_1_status_mxr = io_dpath_status_mxr;
  assign io_requestor_1_status_pum = io_dpath_status_pum;
  assign io_requestor_1_status_mprv = io_dpath_status_mprv;
  assign io_requestor_1_status_xs = io_dpath_status_xs;
  assign io_requestor_1_status_fs = io_dpath_status_fs;
  assign io_requestor_1_status_mpp = io_dpath_status_mpp;
  assign io_requestor_1_status_hpp = io_dpath_status_hpp;
  assign io_requestor_1_status_spp = io_dpath_status_spp;
  assign io_requestor_1_status_mpie = io_dpath_status_mpie;
  assign io_requestor_1_status_hpie = io_dpath_status_hpie;
  assign io_requestor_1_status_spie = io_dpath_status_spie;
  assign io_requestor_1_status_upie = io_dpath_status_upie;
  assign io_requestor_1_status_mie = io_dpath_status_mie;
  assign io_requestor_1_status_hie = io_dpath_status_hie;
  assign io_requestor_1_status_sie = io_dpath_status_sie;
  assign io_requestor_1_status_uie = io_dpath_status_uie;
  assign io_mem_req_valid = T_2580;
  assign io_mem_req_bits_addr = pte_addr[39:0];
  assign io_mem_req_bits_tag = GEN_49;
  assign io_mem_req_bits_cmd = T_2583;
  assign io_mem_req_bits_typ = 3'h3;
  assign io_mem_req_bits_phys = 1'h1;
  assign io_mem_req_bits_data = GEN_123;
  assign io_mem_s1_kill = s1_kill;
  assign io_mem_s1_data = T_2594;
  assign io_mem_invalidate_lr = 1'h0;
  assign T_2207 = r_req_addr[26:18];
  assign T_2208 = r_req_addr[26:9];
  assign vpn_idxs_1 = T_2208[8:0];
  assign vpn_idxs_2 = r_req_addr[8:0];
  assign T_2211 = count & 2'h1;
  assign T_2213 = count >= 2'h2;
  assign T_2217 = T_2211 >= 2'h1;
  assign T_2218 = T_2217 ? vpn_idxs_1 : T_2207;
  assign vpn_idx = T_2213 ? vpn_idxs_2 : T_2218;
  assign arb_clock = clock;
  assign arb_reset = reset;
  assign arb_io_in_0_valid = io_requestor_0_req_valid;
  assign arb_io_in_0_bits_prv = io_requestor_0_req_bits_prv;
  assign arb_io_in_0_bits_pum = io_requestor_0_req_bits_pum;
  assign arb_io_in_0_bits_mxr = io_requestor_0_req_bits_mxr;
  assign arb_io_in_0_bits_addr = io_requestor_0_req_bits_addr;
  assign arb_io_in_0_bits_store = io_requestor_0_req_bits_store;
  assign arb_io_in_0_bits_fetch = io_requestor_0_req_bits_fetch;
  assign arb_io_in_1_valid = io_requestor_1_req_valid;
  assign arb_io_in_1_bits_prv = io_requestor_1_req_bits_prv;
  assign arb_io_in_1_bits_pum = io_requestor_1_req_bits_pum;
  assign arb_io_in_1_bits_mxr = io_requestor_1_req_bits_mxr;
  assign arb_io_in_1_bits_addr = io_requestor_1_req_bits_addr;
  assign arb_io_in_1_bits_store = io_requestor_1_req_bits_store;
  assign arb_io_in_1_bits_fetch = io_requestor_1_req_bits_fetch;
  assign arb_io_out_ready = T_2226;
  assign T_2226 = state == 3'h0;
  assign T_2251_reserved_for_hardware = T_2273;
  assign T_2251_ppn = T_2272;
  assign T_2251_reserved_for_software = T_2271;
  assign T_2251_d = T_2270;
  assign T_2251_a = T_2269;
  assign T_2251_g = T_2268;
  assign T_2251_u = T_2267;
  assign T_2251_x = T_2266;
  assign T_2251_w = T_2265;
  assign T_2251_r = T_2264;
  assign T_2251_v = T_2263;
  assign T_2263 = io_mem_resp_bits_data[0];
  assign T_2264 = io_mem_resp_bits_data[1];
  assign T_2265 = io_mem_resp_bits_data[2];
  assign T_2266 = io_mem_resp_bits_data[3];
  assign T_2267 = io_mem_resp_bits_data[4];
  assign T_2268 = io_mem_resp_bits_data[5];
  assign T_2269 = io_mem_resp_bits_data[6];
  assign T_2270 = io_mem_resp_bits_data[7];
  assign T_2271 = io_mem_resp_bits_data[9:8];
  assign T_2272 = io_mem_resp_bits_data[47:10];
  assign T_2273 = io_mem_resp_bits_data[63:48];
  assign T_2298_reserved_for_hardware = T_2273;
  assign T_2298_ppn = T_2272;
  assign T_2298_reserved_for_software = T_2271;
  assign T_2298_d = T_2270;
  assign T_2298_a = T_2269;
  assign T_2298_g = T_2268;
  assign T_2298_u = T_2267;
  assign T_2298_x = T_2266;
  assign T_2298_w = T_2265;
  assign T_2298_r = T_2264;
  assign T_2298_v = T_2263;
  assign pte_reserved_for_hardware = T_2298_reserved_for_hardware;
  assign pte_ppn = {{18'd0}, T_2332};
  assign pte_reserved_for_software = T_2298_reserved_for_software;
  assign pte_d = T_2298_d;
  assign pte_a = T_2298_a;
  assign pte_g = T_2298_g;
  assign pte_u = T_2298_u;
  assign pte_x = T_2298_x;
  assign pte_w = T_2298_w;
  assign pte_r = T_2298_r;
  assign pte_v = GEN_2;
  assign T_2332 = T_2251_ppn[19:0];
  assign T_2333 = T_2251_ppn[37:20];
  assign T_2335 = T_2333 != 18'h0;
  assign GEN_2 = T_2335 ? 1'h0 : T_2298_v;
  assign T_2337 = {r_pte_ppn,vpn_idx};
  assign GEN_113 = {{3'd0}, T_2337};
  assign pte_addr = GEN_113 << 3;
  assign T_2338 = arb_io_out_ready & arb_io_out_valid;
  assign GEN_3 = T_2338 ? arb_io_out_bits_prv : r_req_prv;
  assign GEN_4 = T_2338 ? arb_io_out_bits_pum : r_req_pum;
  assign GEN_5 = T_2338 ? arb_io_out_bits_mxr : r_req_mxr;
  assign GEN_6 = T_2338 ? arb_io_out_bits_addr : r_req_addr;
  assign GEN_7 = T_2338 ? arb_io_out_bits_store : r_req_store;
  assign GEN_8 = T_2338 ? arb_io_out_bits_fetch : r_req_fetch;
  assign GEN_9 = T_2338 ? arb_io_chosen : r_req_dest;
  assign GEN_10 = T_2338 ? io_dpath_ptbr_ppn : r_pte_ppn;
  assign GEN_114 = {{18'd0}, T_2349_0};
  assign T_2359 = GEN_114 == pte_addr;
  assign GEN_115 = {{18'd0}, T_2349_1};
  assign T_2360 = GEN_115 == pte_addr;
  assign GEN_116 = {{18'd0}, T_2349_2};
  assign T_2361 = GEN_116 == pte_addr;
  assign GEN_117 = {{18'd0}, T_2349_3};
  assign T_2362 = GEN_117 == pte_addr;
  assign GEN_118 = {{18'd0}, T_2349_4};
  assign T_2363 = GEN_118 == pte_addr;
  assign GEN_119 = {{18'd0}, T_2349_5};
  assign T_2364 = GEN_119 == pte_addr;
  assign GEN_120 = {{18'd0}, T_2349_6};
  assign T_2365 = GEN_120 == pte_addr;
  assign GEN_121 = {{18'd0}, T_2349_7};
  assign T_2366 = GEN_121 == pte_addr;
  assign T_2367 = {T_2360,T_2359};
  assign T_2368 = {T_2362,T_2361};
  assign T_2369 = {T_2368,T_2367};
  assign T_2370 = {T_2364,T_2363};
  assign T_2371 = {T_2366,T_2365};
  assign T_2372 = {T_2371,T_2370};
  assign T_2373 = {T_2372,T_2369};
  assign T_2374 = T_2373 & T_2342;
  assign T_2376 = T_2374 != 8'h0;
  assign T_2378 = pte_r == 1'h0;
  assign T_2379 = pte_v & T_2378;
  assign T_2381 = pte_w == 1'h0;
  assign T_2382 = T_2379 & T_2381;
  assign T_2384 = pte_x == 1'h0;
  assign T_2385 = T_2382 & T_2384;
  assign T_2386 = io_mem_resp_valid & T_2385;
  assign T_2388 = T_2376 == 1'h0;
  assign T_2389 = T_2386 & T_2388;
  assign T_2390 = ~ T_2342;
  assign T_2392 = T_2390 == 8'h0;
  assign T_2394 = T_2340 >> 1'h1;
  assign T_2395 = T_2394[0];
  assign T_2396 = {1'h1,T_2395};
  assign T_2397 = T_2340 >> T_2396;
  assign T_2398 = T_2397[0];
  assign T_2399 = {T_2396,T_2398};
  assign T_2400 = T_2340 >> T_2399;
  assign T_2401 = T_2400[0];
  assign T_2402 = {T_2399,T_2401};
  assign T_2403 = T_2402[2:0];
  assign T_2405 = T_2390[0];
  assign T_2406 = T_2390[1];
  assign T_2407 = T_2390[2];
  assign T_2408 = T_2390[3];
  assign T_2409 = T_2390[4];
  assign T_2410 = T_2390[5];
  assign T_2411 = T_2390[6];
  assign T_2421 = T_2411 ? 3'h6 : 3'h7;
  assign T_2422 = T_2410 ? 3'h5 : T_2421;
  assign T_2423 = T_2409 ? 3'h4 : T_2422;
  assign T_2424 = T_2408 ? 3'h3 : T_2423;
  assign T_2425 = T_2407 ? 3'h2 : T_2424;
  assign T_2426 = T_2406 ? 3'h1 : T_2425;
  assign T_2427 = T_2405 ? 3'h0 : T_2426;
  assign T_2428 = T_2392 ? T_2403 : T_2427;
  assign T_2430 = 8'h1 << T_2428;
  assign T_2431 = T_2342 | T_2430;
  assign GEN_0 = pte_addr[31:0];
  assign GEN_11 = 3'h0 == T_2428 ? GEN_0 : T_2349_0;
  assign GEN_12 = 3'h1 == T_2428 ? GEN_0 : T_2349_1;
  assign GEN_13 = 3'h2 == T_2428 ? GEN_0 : T_2349_2;
  assign GEN_14 = 3'h3 == T_2428 ? GEN_0 : T_2349_3;
  assign GEN_15 = 3'h4 == T_2428 ? GEN_0 : T_2349_4;
  assign GEN_16 = 3'h5 == T_2428 ? GEN_0 : T_2349_5;
  assign GEN_17 = 3'h6 == T_2428 ? GEN_0 : T_2349_6;
  assign GEN_18 = 3'h7 == T_2428 ? GEN_0 : T_2349_7;
  assign GEN_1 = pte_ppn[19:0];
  assign GEN_19 = 3'h0 == T_2428 ? GEN_1 : T_2357_0;
  assign GEN_20 = 3'h1 == T_2428 ? GEN_1 : T_2357_1;
  assign GEN_21 = 3'h2 == T_2428 ? GEN_1 : T_2357_2;
  assign GEN_22 = 3'h3 == T_2428 ? GEN_1 : T_2357_3;
  assign GEN_23 = 3'h4 == T_2428 ? GEN_1 : T_2357_4;
  assign GEN_24 = 3'h5 == T_2428 ? GEN_1 : T_2357_5;
  assign GEN_25 = 3'h6 == T_2428 ? GEN_1 : T_2357_6;
  assign GEN_26 = 3'h7 == T_2428 ? GEN_1 : T_2357_7;
  assign GEN_27 = T_2389 ? T_2431 : T_2342;
  assign GEN_28 = T_2389 ? GEN_11 : T_2349_0;
  assign GEN_29 = T_2389 ? GEN_12 : T_2349_1;
  assign GEN_30 = T_2389 ? GEN_13 : T_2349_2;
  assign GEN_31 = T_2389 ? GEN_14 : T_2349_3;
  assign GEN_32 = T_2389 ? GEN_15 : T_2349_4;
  assign GEN_33 = T_2389 ? GEN_16 : T_2349_5;
  assign GEN_34 = T_2389 ? GEN_17 : T_2349_6;
  assign GEN_35 = T_2389 ? GEN_18 : T_2349_7;
  assign GEN_36 = T_2389 ? GEN_19 : T_2357_0;
  assign GEN_37 = T_2389 ? GEN_20 : T_2357_1;
  assign GEN_38 = T_2389 ? GEN_21 : T_2357_2;
  assign GEN_39 = T_2389 ? GEN_22 : T_2357_3;
  assign GEN_40 = T_2389 ? GEN_23 : T_2357_4;
  assign GEN_41 = T_2389 ? GEN_24 : T_2357_5;
  assign GEN_42 = T_2389 ? GEN_25 : T_2357_6;
  assign GEN_43 = T_2389 ? GEN_26 : T_2357_7;
  assign T_2432 = state == 3'h1;
  assign T_2433 = T_2376 & T_2432;
  assign T_2434 = T_2374[7:4];
  assign T_2435 = T_2374[3:0];
  assign T_2437 = T_2434 != 4'h0;
  assign T_2438 = T_2434 | T_2435;
  assign T_2439 = T_2438[3:2];
  assign T_2440 = T_2438[1:0];
  assign T_2442 = T_2439 != 2'h0;
  assign T_2443 = T_2439 | T_2440;
  assign T_2444 = T_2443[1];
  assign T_2445 = {T_2442,T_2444};
  assign T_2446 = {T_2437,T_2445};
  assign T_2448 = T_2446[2];
  assign T_2450 = T_2448 == 1'h0;
  assign T_2452 = 2'h1 << 1'h1;
  assign GEN_122 = {{6'd0}, T_2452};
  assign T_2453 = T_2340 | GEN_122;
  assign T_2454 = ~ T_2340;
  assign T_2455 = T_2454 | GEN_122;
  assign T_2456 = ~ T_2455;
  assign T_2457 = T_2450 ? T_2453 : T_2456;
  assign T_2458 = {1'h1,T_2448};
  assign T_2459 = T_2446[1];
  assign T_2461 = T_2459 == 1'h0;
  assign T_2463 = 4'h1 << T_2458;
  assign GEN_124 = {{4'd0}, T_2463};
  assign T_2464 = T_2457 | GEN_124;
  assign T_2465 = ~ T_2457;
  assign T_2466 = T_2465 | GEN_124;
  assign T_2467 = ~ T_2466;
  assign T_2468 = T_2461 ? T_2464 : T_2467;
  assign T_2469 = {T_2458,T_2459};
  assign T_2470 = T_2446[0];
  assign T_2472 = T_2470 == 1'h0;
  assign T_2474 = 8'h1 << T_2469;
  assign T_2475 = T_2468 | T_2474;
  assign T_2476 = ~ T_2468;
  assign T_2477 = T_2476 | T_2474;
  assign T_2478 = ~ T_2477;
  assign T_2479 = T_2472 ? T_2475 : T_2478;
  assign GEN_44 = T_2433 ? T_2479 : T_2340;
  assign GEN_45 = io_dpath_invalidate ? 8'h0 : GEN_27;
  assign T_2483 = count < 2'h2;
  assign pte_cache_hit = T_2376 & T_2483;
  assign T_2484 = T_2374[0];
  assign T_2485 = T_2374[1];
  assign T_2486 = T_2374[2];
  assign T_2487 = T_2374[3];
  assign T_2488 = T_2374[4];
  assign T_2489 = T_2374[5];
  assign T_2490 = T_2374[6];
  assign T_2491 = T_2374[7];
  assign T_2493 = T_2484 ? T_2357_0 : 20'h0;
  assign T_2495 = T_2485 ? T_2357_1 : 20'h0;
  assign T_2497 = T_2486 ? T_2357_2 : 20'h0;
  assign T_2499 = T_2487 ? T_2357_3 : 20'h0;
  assign T_2501 = T_2488 ? T_2357_4 : 20'h0;
  assign T_2503 = T_2489 ? T_2357_5 : 20'h0;
  assign T_2505 = T_2490 ? T_2357_6 : 20'h0;
  assign T_2507 = T_2491 ? T_2357_7 : 20'h0;
  assign T_2509 = T_2493 | T_2495;
  assign T_2510 = T_2509 | T_2497;
  assign T_2511 = T_2510 | T_2499;
  assign T_2512 = T_2511 | T_2501;
  assign T_2513 = T_2512 | T_2503;
  assign T_2514 = T_2513 | T_2505;
  assign T_2515 = T_2514 | T_2507;
  assign pte_cache_data = T_2515;
  assign T_2541_reserved_for_hardware = T_2565;
  assign T_2541_ppn = T_2564;
  assign T_2541_reserved_for_software = T_2563;
  assign T_2541_d = T_2562;
  assign T_2541_a = T_2561;
  assign T_2541_g = T_2560;
  assign T_2541_u = T_2559;
  assign T_2541_x = T_2558;
  assign T_2541_w = T_2557;
  assign T_2541_r = T_2556;
  assign T_2541_v = T_2555;
  assign T_2554 = 64'h0;
  assign T_2555 = T_2554[0];
  assign T_2556 = T_2554[1];
  assign T_2557 = T_2554[2];
  assign T_2558 = T_2554[3];
  assign T_2559 = T_2554[4];
  assign T_2560 = T_2554[5];
  assign T_2561 = T_2554[6];
  assign T_2562 = T_2554[7];
  assign T_2563 = T_2554[9:8];
  assign T_2564 = T_2554[47:10];
  assign T_2565 = T_2554[63:48];
  assign pte_wdata_reserved_for_hardware = T_2541_reserved_for_hardware;
  assign pte_wdata_ppn = T_2541_ppn;
  assign pte_wdata_reserved_for_software = T_2541_reserved_for_software;
  assign pte_wdata_d = r_req_store;
  assign pte_wdata_a = 1'h1;
  assign pte_wdata_g = T_2541_g;
  assign pte_wdata_u = T_2541_u;
  assign pte_wdata_x = T_2541_x;
  assign pte_wdata_w = T_2541_w;
  assign pte_wdata_r = T_2541_r;
  assign pte_wdata_v = T_2541_v;
  assign T_2579 = state == 3'h4;
  assign T_2580 = T_2432 | T_2579;
  assign T_2583 = T_2579 ? 5'ha : 5'h0;
  assign T_2585 = {pte_wdata_r,pte_wdata_v};
  assign T_2586 = {pte_wdata_u,pte_wdata_x};
  assign T_2587 = {T_2586,pte_wdata_w};
  assign T_2588 = {T_2587,T_2585};
  assign T_2589 = {pte_wdata_d,pte_wdata_a};
  assign T_2590 = {T_2589,pte_wdata_g};
  assign T_2591 = {pte_wdata_reserved_for_hardware,pte_wdata_ppn};
  assign T_2592 = {T_2591,pte_wdata_reserved_for_software};
  assign T_2593 = {T_2592,T_2590};
  assign T_2594 = {T_2593,T_2588};
  assign T_2596 = pte_addr[49:30];
  assign T_2597 = r_req_addr[17:0];
  assign resp_ppns_0 = {T_2596,T_2597};
  assign T_2598 = pte_addr[49:21];
  assign resp_ppns_1 = {T_2598,vpn_idxs_2};
  assign resp_ppns_2 = pte_addr[49:12];
  assign T_2600 = state == 3'h7;
  assign T_2602 = r_req_dest == 1'h0;
  assign T_2603 = T_2600 & T_2602;
  assign T_2612 = T_2217 ? resp_ppns_1 : resp_ppns_0;
  assign T_2613 = T_2213 ? resp_ppns_2 : T_2612;
  assign T_2617 = T_2600 & r_req_dest;
  assign T_2628 = 3'h0 == state;
  assign GEN_46 = arb_io_out_valid ? 3'h1 : state;
  assign GEN_47 = T_2628 ? GEN_46 : state;
  assign GEN_48 = T_2628 ? 2'h0 : count;
  assign T_2630 = 3'h1 == state;
  assign T_2633 = count + 2'h1;
  assign T_2634 = T_2633[1:0];
  assign GEN_50 = pte_cache_hit ? 3'h1 : GEN_47;
  assign GEN_51 = pte_cache_hit ? T_2634 : GEN_48;
  assign GEN_52 = pte_cache_hit ? {{18'd0}, pte_cache_data} : GEN_10;
  assign T_2636 = pte_cache_hit == 1'h0;
  assign T_2637 = T_2636 & io_mem_req_ready;
  assign GEN_53 = T_2637 ? 3'h2 : GEN_50;
  assign GEN_54 = T_2630 ? pte_cache_hit : 1'h0;
  assign GEN_55 = T_2630 ? GEN_53 : GEN_47;
  assign GEN_56 = T_2630 ? GEN_51 : GEN_48;
  assign GEN_57 = T_2630 ? GEN_52 : GEN_10;
  assign T_2638 = 3'h2 == state;
  assign GEN_58 = io_mem_xcpt_pf_ld ? 1'h0 : r_pte_v;
  assign GEN_59 = io_mem_xcpt_pf_ld ? 3'h7 : 3'h3;
  assign GEN_60 = T_2638 ? GEN_59 : GEN_55;
  assign GEN_61 = T_2638 ? GEN_58 : r_pte_v;
  assign T_2640 = 3'h3 == state;
  assign GEN_62 = io_mem_s2_nack ? 3'h1 : GEN_60;
  assign T_2641 = pte_x & r_req_mxr;
  assign T_2642 = pte_r | T_2641;
  assign T_2643 = r_req_store ? pte_w : T_2642;
  assign T_2644 = r_req_fetch ? pte_x : T_2643;
  assign T_2646 = r_req_pum == 1'h0;
  assign T_2647 = r_req_prv[0];
  assign T_2648 = pte_u ? T_2646 : T_2647;
  assign T_2651 = pte_x & T_2381;
  assign T_2652 = pte_r | T_2651;
  assign T_2653 = pte_v & T_2652;
  assign T_2654 = T_2653 & T_2648;
  assign T_2655 = T_2654 & T_2644;
  assign T_2657 = pte_a == 1'h0;
  assign T_2659 = pte_d == 1'h0;
  assign T_2660 = r_req_store & T_2659;
  assign T_2661 = T_2657 | T_2660;
  assign T_2662 = T_2655 & T_2661;
  assign GEN_63 = T_2662 ? 3'h4 : 3'h7;
  assign T_2664 = T_2662 == 1'h0;
  assign GEN_64 = T_2664 ? pte_reserved_for_hardware : r_pte_reserved_for_hardware;
  assign GEN_65 = T_2664 ? pte_ppn : GEN_57;
  assign GEN_66 = T_2664 ? pte_reserved_for_software : r_pte_reserved_for_software;
  assign GEN_67 = T_2664 ? pte_d : r_pte_d;
  assign GEN_68 = T_2664 ? pte_a : r_pte_a;
  assign GEN_69 = T_2664 ? pte_g : r_pte_g;
  assign GEN_70 = T_2664 ? pte_u : r_pte_u;
  assign GEN_71 = T_2664 ? pte_x : r_pte_x;
  assign GEN_72 = T_2664 ? pte_w : r_pte_w;
  assign GEN_73 = T_2664 ? pte_r : r_pte_r;
  assign GEN_74 = T_2664 ? pte_v : GEN_61;
  assign T_2676 = T_2385 & T_2483;
  assign GEN_75 = T_2676 ? 3'h1 : GEN_63;
  assign GEN_76 = T_2676 ? T_2634 : GEN_56;
  assign GEN_77 = io_mem_resp_valid ? GEN_75 : GEN_62;
  assign GEN_78 = io_mem_resp_valid ? GEN_64 : r_pte_reserved_for_hardware;
  assign GEN_79 = io_mem_resp_valid ? GEN_65 : GEN_57;
  assign GEN_80 = io_mem_resp_valid ? GEN_66 : r_pte_reserved_for_software;
  assign GEN_81 = io_mem_resp_valid ? GEN_67 : r_pte_d;
  assign GEN_82 = io_mem_resp_valid ? GEN_68 : r_pte_a;
  assign GEN_83 = io_mem_resp_valid ? GEN_69 : r_pte_g;
  assign GEN_84 = io_mem_resp_valid ? GEN_70 : r_pte_u;
  assign GEN_85 = io_mem_resp_valid ? GEN_71 : r_pte_x;
  assign GEN_86 = io_mem_resp_valid ? GEN_72 : r_pte_w;
  assign GEN_87 = io_mem_resp_valid ? GEN_73 : r_pte_r;
  assign GEN_88 = io_mem_resp_valid ? GEN_74 : GEN_61;
  assign GEN_89 = io_mem_resp_valid ? GEN_76 : GEN_56;
  assign GEN_90 = T_2640 ? GEN_77 : GEN_60;
  assign GEN_91 = T_2640 ? GEN_78 : r_pte_reserved_for_hardware;
  assign GEN_92 = T_2640 ? GEN_79 : GEN_57;
  assign GEN_93 = T_2640 ? GEN_80 : r_pte_reserved_for_software;
  assign GEN_94 = T_2640 ? GEN_81 : r_pte_d;
  assign GEN_95 = T_2640 ? GEN_82 : r_pte_a;
  assign GEN_96 = T_2640 ? GEN_83 : r_pte_g;
  assign GEN_97 = T_2640 ? GEN_84 : r_pte_u;
  assign GEN_98 = T_2640 ? GEN_85 : r_pte_x;
  assign GEN_99 = T_2640 ? GEN_86 : r_pte_w;
  assign GEN_100 = T_2640 ? GEN_87 : r_pte_r;
  assign GEN_101 = T_2640 ? GEN_88 : GEN_61;
  assign GEN_102 = T_2640 ? GEN_89 : GEN_56;
  assign T_2680 = 3'h4 == state;
  assign GEN_103 = io_mem_req_ready ? 3'h5 : GEN_90;
  assign GEN_104 = T_2680 ? GEN_103 : GEN_90;
  assign T_2681 = 3'h5 == state;
  assign GEN_105 = io_mem_xcpt_pf_st ? 1'h0 : GEN_101;
  assign GEN_106 = io_mem_xcpt_pf_st ? 3'h7 : 3'h6;
  assign GEN_107 = T_2681 ? GEN_106 : GEN_104;
  assign GEN_108 = T_2681 ? GEN_105 : GEN_101;
  assign T_2683 = 3'h6 == state;
  assign GEN_109 = io_mem_s2_nack ? 3'h4 : GEN_107;
  assign GEN_110 = io_mem_resp_valid ? 3'h1 : GEN_109;
  assign GEN_111 = T_2683 ? GEN_110 : GEN_107;
  assign T_2684 = 3'h7 == state;
  assign GEN_112 = T_2684 ? 3'h0 : GEN_111;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_125 = {1{$random}};
  state = GEN_125[2:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_126 = {1{$random}};
  count = GEN_126[1:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_127 = {1{$random}};
  s1_kill = GEN_127[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_128 = {1{$random}};
  r_req_prv = GEN_128[1:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_129 = {1{$random}};
  r_req_pum = GEN_129[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_130 = {1{$random}};
  r_req_mxr = GEN_130[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_131 = {1{$random}};
  r_req_addr = GEN_131[26:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_132 = {1{$random}};
  r_req_store = GEN_132[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_133 = {1{$random}};
  r_req_fetch = GEN_133[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_134 = {1{$random}};
  r_req_dest = GEN_134[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_135 = {1{$random}};
  r_pte_reserved_for_hardware = GEN_135[15:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_136 = {2{$random}};
  r_pte_ppn = GEN_136[37:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_137 = {1{$random}};
  r_pte_reserved_for_software = GEN_137[1:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_138 = {1{$random}};
  r_pte_d = GEN_138[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_139 = {1{$random}};
  r_pte_a = GEN_139[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_140 = {1{$random}};
  r_pte_g = GEN_140[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_141 = {1{$random}};
  r_pte_u = GEN_141[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_142 = {1{$random}};
  r_pte_x = GEN_142[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_143 = {1{$random}};
  r_pte_w = GEN_143[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_144 = {1{$random}};
  r_pte_r = GEN_144[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_145 = {1{$random}};
  r_pte_v = GEN_145[0:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_146 = {1{$random}};
  T_2340 = GEN_146[7:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_147 = {1{$random}};
  T_2342 = GEN_147[7:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_148 = {1{$random}};
  T_2349_0 = GEN_148[31:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_149 = {1{$random}};
  T_2349_1 = GEN_149[31:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_150 = {1{$random}};
  T_2349_2 = GEN_150[31:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_151 = {1{$random}};
  T_2349_3 = GEN_151[31:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_152 = {1{$random}};
  T_2349_4 = GEN_152[31:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_153 = {1{$random}};
  T_2349_5 = GEN_153[31:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_154 = {1{$random}};
  T_2349_6 = GEN_154[31:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_155 = {1{$random}};
  T_2349_7 = GEN_155[31:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_156 = {1{$random}};
  T_2357_0 = GEN_156[19:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_157 = {1{$random}};
  T_2357_1 = GEN_157[19:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_158 = {1{$random}};
  T_2357_2 = GEN_158[19:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_159 = {1{$random}};
  T_2357_3 = GEN_159[19:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_160 = {1{$random}};
  T_2357_4 = GEN_160[19:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_161 = {1{$random}};
  T_2357_5 = GEN_161[19:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_162 = {1{$random}};
  T_2357_6 = GEN_162[19:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_163 = {1{$random}};
  T_2357_7 = GEN_163[19:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_164 = {1{$random}};
  GEN_49 = GEN_164[6:0];
  `endif
  `ifdef RANDOMIZE_REG_INIT
  GEN_165 = {2{$random}};
  GEN_123 = GEN_165[63:0];
  `endif
  end
`endif
  always @(posedge clock) begin
    if(reset) begin
      state <= 3'h0;
    end else begin 
      if(T_2684) begin // state == 7, state == done
        state <= 3'h0; // state <= ready
      end else begin
        if(T_2683) begin // state == 6, state == wait2_dirty
          if(io_mem_resp_valid) begin
            state <= 3'h1; // state <= req
          end else begin
            if(io_mem_s2_nack) begin 
              state <= 3'h4; // state <= set_dirty
            end /*else begin
              if(T_2681) begin // state == 5, state == wait1_dirty
                if(io_mem_xcpt_pf_st) begin
                  state <= 3'h7; // state <= done
                end else begin
                  state <= 3'h6; // state <= wait2_dirty
                end
              end else begin
                if(T_2680) begin // state == 4, state == set_dirty
                  if(io_mem_req_ready) begin
                    state <= 3'h5; // state <= wait1_dirty
                  end else begin
                    if(T_2640) begin // state == 3, state == wait2
                      if(io_mem_resp_valid) begin
                        if(T_2676) begin // count < 2 && (v && !r && !w && !x), 即非叶子页表
                          state <= 3'h1; // state <= req
                        end else begin
                          if(T_2662) begin // access_ok，权限检查
                            state <= 3'h4; // state <= set_dirty
                          end else begin
                            state <= 3'h7; // state <= done
                          end
                        end
                      end else begin
                        if(io_mem_s2_nack) begin
                          state <= 3'h1; // state <= req
                        end else begin
                          if(T_2638) begin // state == 2, state == wait1
                            if(io_mem_xcpt_pf_ld) begin
                              state <= 3'h7;
                            end else begin
                              state <= 3'h3;
                            end
                          end else begin
                            if(T_2630) begin
                              if(T_2637) begin
                                state <= 3'h2;
                              end else begin
                                if(pte_cache_hit) begin
                                  state <= 3'h1;
                                end else begin
                                  if(T_2628) begin
                                    if(arb_io_out_valid) begin
                                      state <= 3'h1;
                                    end
                                  end
                                end
                              end
                            end else begin
                              if(T_2628) begin
                                if(arb_io_out_valid) begin
                                  state <= 3'h1;
                                end
                              end
                            end
                          end
                        end
                      end
                    end else begin
                      if(T_2638) begin // state == 2, state == wait1
                        if(io_mem_xcpt_pf_ld) begin
                          state <= 3'h7; // state <= done
                        end else begin
                          state <= 3'h3; // state <= wait2
                        end
                      end else begin
                        if(T_2630) begin // state == 1, state == req
                          if(T_2637) begin // !pte_cache_hit && io_mem_req_ready
                            state <= 3'h2; // state <= wait1
                          end else begin
                            if(pte_cache_hit) begin 
                              state <= 3'h1; // state <= req
                            end else begin
                              if(T_2628) begin // state == 0, state == ready
                                if(arb_io_out_valid) begin
                                  state <= 3'h1; // state <= req
                                end
                              end
                            end
                          end
                        end else begin
                          if(T_2628) begin // state == 0, state == ready
                            if(arb_io_out_valid) begin
                              state <= 3'h1; // state <= req
                            end
                          end
                        end
                      end
                    end
                  end
                end else begin
                  if(T_2640) begin // state == 
                    if(io_mem_resp_valid) begin
                      if(T_2676) begin
                        state <= 3'h1;
                      end else begin
                        if(T_2662) begin
                          state <= 3'h4;
                        end else begin
                          state <= 3'h7;
                        end
                      end
                    end else begin
                      if(io_mem_s2_nack) begin
                        state <= 3'h1;
                      end else begin
                        if(T_2638) begin
                          if(io_mem_xcpt_pf_ld) begin
                            state <= 3'h7;
                          end else begin
                            state <= 3'h3;
                          end
                        end else begin
                          if(T_2630) begin
                            if(T_2637) begin
                              state <= 3'h2;
                            end else begin
                              if(pte_cache_hit) begin
                                state <= 3'h1;
                              end else begin
                                state <= GEN_47;
                              end
                            end
                          end else begin
                            state <= GEN_47;
                          end
                        end
                      end
                    end
                  end else begin
                    if(T_2638) begin
                      if(io_mem_xcpt_pf_ld) begin
                        state <= 3'h7;
                      end else begin
                        state <= 3'h3;
                      end
                    end else begin
                      if(T_2630) begin
                        if(T_2637) begin
                          state <= 3'h2;
                        end else begin
                          if(pte_cache_hit) begin
                            state <= 3'h1;
                          end else begin
                            state <= GEN_47;
                          end
                        end
                      end else begin
                        state <= GEN_47;
                      end
                    end
                  end
                end
              end
            end*/
          end
        end else begin
          if(T_2681) begin // state == 5, state == wait1_dirty
            if(io_mem_xcpt_pf_st) begin
              state <= 3'h7; // state <= done
            end else begin
              state <= 3'h6; // state <= wait2_dirty
            end
          end else begin
            if(T_2680) begin // state == 4, state == set_dirty
              if(io_mem_req_ready) begin
                state <= 3'h5; // state <= wait1_dirty
              end /*else begin
                if(T_2640) begin // state == 3
                  if(io_mem_resp_valid) begin
                    if(T_2676) begin
                      state <= 3'h1;
                    end else begin
                      if(T_2662) begin
                        state <= 3'h4;
                      end else begin
                        state <= 3'h7;
                      end
                    end
                  end else begin
                    if(io_mem_s2_nack) begin
                      state <= 3'h1;
                    end else begin
                      state <= GEN_60;
                    end
                  end
                end else begin
                  state <= GEN_60;
                end
              end*/
            end else begin
              if(T_2640) begin // state == 3, state == wait2
                if(io_mem_resp_valid) begin
                  if(T_2676) begin // (v && !r && !w && !x) && count < 2, 即非叶子页表
                    state <= 3'h1; // state <= req
                  end else begin
                    if(T_2662) begin // access_ok && (!d && req_store_ || !a)
                      state <= 3'h4; // state <= wait2
                    end else begin
                      state <= 3'h7; // state <= done
                    end
                  end
                end else begin
                  if(io_mem_s2_nack) begin
                    state <= 3'h1; // state <= req
                  end/* else begin
                    state <= GEN_60;
                  end*/
                end
              end else begin // state == 1, state == 0
                state <= GEN_60;
              end
            end
          end
        end
      end
    end


    // set registers' value
    if(1'h0) begin
    end else begin
      if(T_2640) begin // state == 3, state == wait2
        if(io_mem_resp_valid) begin
          if(T_2676) begin // (v && !r && !w && !x) && count < 2, 即非叶子页表
            count <= T_2634; // count ++
          end/* else begin
            if(T_2630) begin // state == 1,
              if(pte_cache_hit) begin
                count <= T_2634; // count ++
              end else begin
                if(T_2628) begin // state == 0, 
                  count <= 2'h0;
                end
              end
            end else begin
              if(T_2628) begin
                count <= 2'h0;
              end
            end
          end
        end else begin
          if(T_2630) begin
            if(pte_cache_hit) begin
              count <= T_2634;
            end else begin
              if(T_2628) begin
                count <= 2'h0;
              end
            end
          end else begin
            if(T_2628) begin
              count <= 2'h0;
            end
          end*/
        end
      end else begin
        if(T_2630) begin // state == 1, state == req
          if(pte_cache_hit) begin
            count <= T_2634; // count++
          end else begin
            count <= GEN_48; // GEN_48 = state == 3'h0 ? 2'h0 : count
          end
        end else begin // state == 0, state == ready
          count <= GEN_48;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_2630) begin // state == 1, state == req
        s1_kill <= pte_cache_hit; 
      end else begin
        s1_kill <= 1'h0; 
      end
    end
    if(1'h0) begin
    end else begin
      if(T_2338) begin // arb_io_out_ready && arb_io_out_valid
        // 缓存请求
        r_req_prv <= arb_io_out_bits_prv;
        r_req_pum <= arb_io_out_bits_pum;
        r_req_mxr <= arb_io_out_bits_mxr;
        r_req_addr <= arb_io_out_bits_addr;
        r_req_store <= arb_io_out_bits_store;
        r_req_fetch <= arb_io_out_bits_fetch;
        r_req_dest <= arb_io_chosen;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_2640) begin // state == 3, state == wait2
        if(io_mem_resp_valid) begin
          if(T_2664) begin // !(access_ok && ((!d && r_req_store) || !a)
            r_pte_reserved_for_hardware <= pte_reserved_for_hardware;
            r_pte_ppn <= pte_ppn;
            r_pte_reserved_for_software <= pte_reserved_for_software;
            r_pte_d <= pte_d;
            r_pte_a <= pte_a;
            r_pte_g <= pte_g;
            r_pte_u <= pte_u;
            r_pte_x <= pte_x;
            r_pte_w <= pte_w;
            r_pte_r <= pte_r;
          end/* else begin
            if(T_2630) begin // state == 1, state == req
              if(pte_cache_hit) begin
                r_pte_ppn <= {{18'd0}, pte_cache_data};
              end else begin
                if(T_2338) begin
                  r_pte_ppn <= io_dpath_ptbr_ppn;
                end
              end
            end else begin
              if(T_2338) begin
                r_pte_ppn <= io_dpath_ptbr_ppn;
              end
            end
          end
        end else begin
          if(T_2630) begin
            if(pte_cache_hit) begin
              r_pte_ppn <= {{18'd0}, pte_cache_data};
            end else begin
              if(T_2338) begin
                r_pte_ppn <= io_dpath_ptbr_ppn;
              end
            end
          end else begin
            if(T_2338) begin
              r_pte_ppn <= io_dpath_ptbr_ppn;
            end
          end*/
        end
      end else begin
        if(T_2630) begin // state == 1, state = req
          if(pte_cache_hit) begin
            r_pte_ppn <= {{18'd0}, pte_cache_data};
          end else begin
            r_pte_ppn <= GEN_10;
          end
        end else begin
          r_pte_ppn <= GEN_10;
        end
      end
    end
    /*
    if(1'h0) begin
    end else begin
      if(T_2640) begin
        if(io_mem_resp_valid) begin
          if(T_2664) begin
            r_pte_reserved_for_hardware <= pte_reserved_for_hardware;
            r_pte_ppn <= pte_ppn;
            r_pte_reserved_for_software <= pte_reserved_for_software;
            r_pte_d <= pte_d;
            r_pte_a <= pte_a;
            r_pte_g <= pte_g;
            r_pte_u <= pte_u;
            r_pte_x <= pte_x;
            r_pte_w <= pte_w;
            r_pte_r <= pte_r;
          end
        end
      end
    end*/
    if(1'h0) begin
    end else begin
      if(T_2681) begin // state == 5, state == wait1_dirty
        if(io_mem_xcpt_pf_st) begin
          r_pte_v <= 1'h0;
        end/* else begin
          if(T_2640) begin // state == 3
            if(io_mem_resp_valid) begin
              if(T_2664) begin
                r_pte_v <= pte_v;
              end else begin
                if(T_2638) begin // state == 2
                  if(io_mem_xcpt_pf_ld) begin
                    r_pte_v <= 1'h0;
                  end
                end
              end
            end else begin
              if(T_2638) begin // state == 2
                if(io_mem_xcpt_pf_ld) begin
                  r_pte_v <= 1'h0;
                end
              end
            end
          end else begin
            if(T_2638) begin // state == 2
              if(io_mem_xcpt_pf_ld) begin
                r_pte_v <= 1'h0;
              end
            end
          end
        end*/
      end else begin
        if(T_2640) begin // state == 3, state == wait2
          if(io_mem_resp_valid) begin
            if(T_2664) begin
              r_pte_v <= pte_v;
            end/* else begin
              if(T_2638) begin // state == 2
                if(io_mem_xcpt_pf_ld) begin
                  r_pte_v <= 1'h0;
                end
              end
            end*/
          end else begin
            r_pte_v <= GEN_61;
          end
        end else begin
          r_pte_v <= GEN_61;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_2433) begin // state == 1 && 缓存命中
        if(T_2472) begin // 
          T_2340 <= T_2475; // 可能是PLRU寄存器
        end else begin
          T_2340 <= T_2478;
        end
      end
    end
    // 设置valid
    if(reset) begin 
      T_2342 <= 8'h0;
    end else begin
      if(io_dpath_invalidate) begin
        T_2342 <= 8'h0;
      end else begin
        if(T_2389) begin // 缓存未命中 && (v & !r & !w & !x) && io_mem_resp_valid
          T_2342 <= T_2431; // 更新valid
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_2389) begin // 缓存未命中 && (v & !r & !w & !x) && io_mem_resp_valid
        // 更新pte_addr, 32位
        if(3'h0 == T_2428) begin
          T_2349_0 <= GEN_0;
        end
        if(3'h1 == T_2428) begin
          T_2349_1 <= GEN_0;
        end
        if(3'h2 == T_2428) begin
          T_2349_2 <= GEN_0;
        end
        if(3'h3 == T_2428) begin
          T_2349_3 <= GEN_0;
        end
        if(3'h4 == T_2428) begin
          T_2349_4 <= GEN_0;
        end
        if(3'h5 == T_2428) begin
          T_2349_5 <= GEN_0;
        end
        if(3'h6 == T_2428) begin
          T_2349_6 <= GEN_0;
        end
        if(3'h7 == T_2428) begin
          T_2349_7 <= GEN_0;
        end
      //////////////////////////////
      // 更新pte_ppn, 20位
        if(3'h0 == T_2428) begin
          T_2357_0 <= GEN_1;
        end
        if(3'h1 == T_2428) begin
          T_2357_1 <= GEN_1;
        end
        if(3'h2 == T_2428) begin
          T_2357_2 <= GEN_1;
        end
        if(3'h3 == T_2428) begin
          T_2357_3 <= GEN_1;
        end
        if(3'h4 == T_2428) begin
          T_2357_4 <= GEN_1;
        end
        if(3'h5 == T_2428) begin
          T_2357_5 <= GEN_1;
        end
        if(3'h6 == T_2428) begin
          T_2357_6 <= GEN_1;
        end
        if(3'h7 == T_2428) begin
          T_2357_7 <= GEN_1;
        end
      end
    end
  end
endmodule